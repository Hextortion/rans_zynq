`timescale 1ns / 1ps
`default_nettype none

`include "rans_if.sv"

package RansTestPackage;
    `include "transaction.sv"
    `include "driver.sv"
endpackage : RansTestPackage